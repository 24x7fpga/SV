class cstrs_challenge;

   // class properties

   // display function
   function void disp();
     
   endfunction // disp

endclass // cstrs_challenge
