class transaction #(parameter N = 4);

   // declare random variables
   // Outputs
    
   // Inputs
  
   // add constraints
  
  
  
   // display function
   function void DISP(string name);
      $display(" %s: <SIGNALS>", name, <SIGNALS>);
   endfunction // DISP

endclass // transaction
