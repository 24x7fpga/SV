class transaction;

   // declare random variables

   // add constraints

   // display function
   function void DISP(string name);
      $display(" %s: < decalre variables>", name, <declare varibles>);
   endfunction // DISP

endclass // transaction
