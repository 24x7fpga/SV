//Interface 

//Declare all the inputs and outputs using logic 
//this may also contain modport and clocking block based on the design

interface intf();
  
  logic a;
  logic b;
  logic c;
  
  logic s;
  logic co;
  
endinterface;
