`include "test.sv"

module tb_diag_zero;
   
   test t1();

endmodule // tb_diag_zero   

