`include "test.sv"

module tb_$ARG;
   
   test t1 ();

endmodule // tb_$ARG   

