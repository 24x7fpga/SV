`include "test.sv"

module tb_non_consecutive;
   
   test t1 ();

endmodule // tb_non_consecutive   

