interface intf();

  //Declare all the inputs and outputs using logic 
  //this may also contain modport and clocking block based on the design

  
endinterface
