interface intf #(parameter int N = 1) (input clk);

   // Outputs
   // Inputs
   
endinterface
